`timescale 1ns / 1ps
`include "defines.vh"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/11/02 14:52:16
// Design Name: 
// Module Name: alu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alu(
	input wire[31:0] a,b,
	input wire[7:0] op,
//	input wire[4:0] sa,
	output reg[31:0] y,
	output reg overflow,
	output wire zero
    );

	wire[31:0] s,bout;
	
	always @(*) begin
		case (op)
			`EXE_AND_OP: y <= a & b; //and
			`EXE_OR_OP: y <= a | b; //or
			`EXE_XOR_OP: y <= a^b; //xor
			`EXE_NOR_OP: y <= ~a^b; //nor
			
			`EXE_ANDI_OP: y <= a & b; //andi
			`EXE_ORI_OP: y <= a | b; //ori
			`EXE_XORI_OP: y <= a^b; //xori
			`EXE_LUI_OP: y <= {b[31:16],{16{1'b0}}}; //lui
			
			default : y <= 32'b0;
		endcase	
	end
	
	assign zero = (y == 32'b0);

	always @(*) begin
		case (op[2:1])
			2'b01:overflow <= a[31] & b[31] & ~s[31] |
							~a[31] & ~b[31] & s[31];
			2'b11:overflow <= ~a[31] & b[31] & s[31] |
							a[31] & ~b[31] & ~s[31];
			default : overflow <= 1'b0;
		endcase	
	end
endmodule

`timescale 1ns / 1ps
`include "defines.vh"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/10/23 15:21:30
// Design Name: 
// Module Name: maindec
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module maindec(
	input wire[5:0] op,
    input wire[5:0] funct,
    input wire[4:0] rt,
	output wire memtoreg,memwrite,
	output wire branch,alusrc,
	output wire regdst,regwrite,
	output wire jump
//	output wire[1:0] aluop
    );
	reg[8:0] controls;
	assign {regwrite,regdst,alusrc,branch,memwrite,memtoreg,jump} = controls;
	always @(*) begin
		case (op)
			//I-TYPE
			`EXE_ANDI:controls <= 7'b1010000;
			`EXE_XORI:controls <= 7'b1010000;
			`EXE_LUI:controls <= 7'b1010000;
			`EXE_ORI:controls <= 7'b1010000; //�������߼�����ָ��
	        
	        `EXE_ADDI:controls <= 7'b1010000;
	        `EXE_ADDIU:controls <= 7'b1010000;
	        `EXE_SLTI:controls <= 7'b1010000;
	        `EXE_SLTIU:controls <= 7'b1010000; // ����������ָ��
	        
	        //R-TYRE
	        `EXE_ADD:controls <= 7'b1100000;
	        `EXE_ADDU:controls <= 7'b1100000;
	        `EXE_SUB:controls <= 7'b1100000;
	        `EXE_SUBU:controls <= 7'b1100000;
	        `EXE_SLT:controls <= 7'b1100000;
	        `EXE_SLTU:controls <= 7'b1100000; //R������ָ��


			6'b100011:controls <= 7'b1010010;//LW
			6'b101011:controls <= 7'b0010100;//SW
			6'b000100:controls <= 7'b0001000;//BEQ
			
			6'b000010:controls <= 7'b0000001;//J
			default:  controls <= 7'b0000000;//illegal op
		endcase
	end
endmodule
